module Minilab1 (
    input wire clk,
    input wire reset_n
);

//8 MACS



//9 FIFOS



endmodule;